/home/alex/FPGALAB/Lab1/lab1/lab1.srcs/sources_1/new/top.sv